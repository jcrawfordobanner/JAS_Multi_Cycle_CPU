module concatinate(
  input notconcatinated,
  output concatinated
);
 assign extended = {4'b0,in,2'b0};
 endmodule
